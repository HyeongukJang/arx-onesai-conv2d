
`define USE_SRAM
`define SRAM_HEX_SIZE 8
`define CRM_HEX_SIZE 0
`define USE_DRAM
`define DRAM_HEX_SIZE 36176
`define HEX_SIZE 36176